//=====================================================
// Project     : SPI (Serial Peripheral Interface)
// File        : sequencer.sv
// Author      : Brahma Ganesh Katrapalli
// Created On  : 18-12-2025
// Revision    : 1.0
// Description : Sequencer controlling transaction flow to driver
//=====================================================

class spi_sequencer extends uvm_sequencer#(spi_transaction);
    `uvm_component_utils(spi_sequencer)
    
    function new(string name="spi_sequencer", uvm_component parent=null);
        super.new(name,parent);
    endfunction

endclass
